module crm();
endmodule
