module clk_reg_div();
endmodule
