module tb();
endmodule
