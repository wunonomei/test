module testcase();
endmodule
